module hassclient



